//design file 
module _4_1mux(input [1:0]a,b,c,d,input s0,s1,output reg[1:0] y);
  always@(*)
    begin
      case({s1,s0})
      2'b00 :y=a;
      2'b01 :y=b;
      2'b10:y=c;
      2'b11:y=d;
        default:y=0;
    endcase
  end
      
endmodule

//test bench file 
module _4_1mux_tb;
  reg [1:0]a,b,c,d;
  reg s0,s1;
  wire [1:0]y;
  _4_1mux uut(a,b,c,d,s0,s1,y);
  initial 
    begin 
      $monitor("time=%0t s0=%b s1=%b y=%b",$time,s0,s1,y);
      a=2'b0;b=2'b1;c=2'b10;d=2'b11;
      #3 s1=1;s0=1;
       #3 s1=0;s0=1;
       #3 s1=0;s0=0;
      #20$finish;
    end
endmodule 
